package CIMulator_PKG;

localparam CIM_ADDRESS_DEPTH = 512;
localparam CIM_ADDR_WIDTH = 8;
localparam CIM_ADDR_AV_WIDTH = CIM_ADDR_WIDTH + 1;

endpackage